class coverfloat_coverage; import coverfloat_pkg::*;

    // constructor (initializes covergroups)
    
    // covergroups and sample functions (probably `include 'd)

endclass