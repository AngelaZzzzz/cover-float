        // all conversion operations
        bins op_cfi    = {[OP_CFI  : OP_CFI  | 32'hF]};
        bins op_fcvtw  = {OP_FCVTW};
        bins op_fcvtwu = {OP_FCVTWU};
        bins op_fcvtl  = {OP_FCVTL};
        bins op_fcvtlu = {OP_FCVTLU};
        bins op_cff    = {[OP_CFF   : OP_CFF   | 32'hF]}; 